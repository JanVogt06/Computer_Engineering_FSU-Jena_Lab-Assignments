/**
 * 4-bit ripple-carry adder.
 *
 * @param i_a input A.
 * @param i_b input B.
 * @param i_carry_in carry in.
 * @param o_s sum.
 * @param o_carry_out carry out.
 **/
module ripple_carry_adder_4 (
    input  logic [3:0] i_a,
    i_b,
    input  logic       i_carry_in,
    output logic [3:0] o_s,
    output logic       o_carry_out
);
    // TODO: implement 4-bit ripple-carry adder
endmodule

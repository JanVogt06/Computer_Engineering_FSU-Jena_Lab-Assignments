/**
 * Gate-level implementation of a full adder.
 *
 * @param i_a input A.
 * @param i_b input B.
 * @param i_carry_in carry in.
 * @param o_s sum.
 * @param o_carry_out carry out.
 **/
module full_adder(
        input  wire i_a,
                    i_b,
                    i_carry_in,
        output wire o_s,
                    o_carry_out
    );

    
endmodule